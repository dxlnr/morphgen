module cpu
endmodule
